//////////////////////////////////////////////////
// Title:   in_hdlc
// Author:
// Date:
//////////////////////////////////////////////////

interface in_hdlc ();
  //Tb
  int ErrCntAssertions;

  //Clock and reset
  logic              Clk;
  logic              Rst;

  // Address
  logic        [2:0] Address;
  logic              WriteEnable;
  logic              ReadEnable;
  logic        [7:0] DataIn;
  logic        [7:0] DataOut;

  // TX
  logic              Tx;
  logic              TxEN;
  logic              Tx_Done;

  // RX
  logic              Rx;
  logic              RxEN;
  logic              Rx_Ready;

  // Tx - internal
  logic             Tx_DataAvail;
  logic             Tx_Full;
  logic       [7:0] Tx_Data;
  logic             Tx_NewByte;
  logic       [7:0] Tx_FrameSize;
  logic             Tx_Enable;
  logic             Tx_AbortedTrans;
  logic             Tx_AbortFrame;
  logic             Tx_ValidFrame;
  logic             Tx_WriteFCS;
  logic             Tx_FCSDone;
  // Rx - internal
  logic       Rx_FlagDetect;
  logic       Rx_Drop;
  logic       Rx_AbortSignal;
  logic       Rx_ValidFrame;
  logic       Rx_FrameError;
  logic       [7:0] Rx_Data;
  logic       Rx_EoF;
  logic       Rx_Overflow;



endinterface
