//////////////////////////////////////////////////
// Title:   testPr_hdlc
// Author:
// Date:
//////////////////////////////////////////////////


program testPr_hdlc(
  in_hdlc uin_hdlc
);

// class data_hdlc;
//   rand logic [0:7] inputValue;
//
//   task get(ref logic [0:7] inputValue);
//     inputValue = inputValue;
//   endtask
// endclass: data_hdlc;
  int TbErrorCnt;
  parameter TX_SC   = 3'b000;
  parameter TX_BUFF = 3'b001;
  parameter RX_SC   = 3'b010;
  parameter RX_BUFF = 3'b011;
  parameter RX_LEN  = 3'b100;

  parameter TX_DONE         = 8'b0000_0001;
  parameter TX_ENABLE       = 8'b0000_0010;
  parameter TX_ABORTFRAME   = 8'b0000_0100;
  parameter TX_ABORTEDTRANS = 8'b0000_1000;
  parameter TX_FULL         = 8'b0001_0000;

  parameter RX_READY        = 8'b0000_0001;
  parameter RX_DROP         = 8'b0000_0010;
  parameter RX_FRAMEERROR   = 8'b0000_0100;
  parameter RX_ABORTSIGNAL  = 8'b0000_1000;
  parameter RX_OVERFLOW     = 8'b0001_0000;
  parameter RX_FCSEN        = 8'b0010_0000;

  int num_loops = 50;



  initial begin
    $display("*************************************************************");
    $display("%t - Starting Test Program", $time);
    $display("*************************************************************");

    init();

    //Tests:
    //Receive();
    //Verification1_Drop();
    //Verification1_Abort();
    //Verification1_Error();
    //Verification17();
    //Verification9();
    //Verification6();
//    Verification8();
    for(int loop = 0; loop < num_loops; loop++) begin
        $display("Random test %d", loop+1);
        random_input();
    end
    $display("*************************************************************");
    $display("%t - Finishing Test Program", $time);
    $display("*************************************************************");
    $stop;
  end

  final begin

    $display("*********************************");
    $display("*                               *");
    $display("* \tAssertion Errors: %0d\t  *", TbErrorCnt + uin_hdlc.ErrCntAssertions);
    $display("*                               *");
    $display("*********************************");

  end

  task init();
    uin_hdlc.Clk         =   1'b0;
    uin_hdlc.Rst         =   1'b0;
    uin_hdlc.Rx          =   1'b0;
    uin_hdlc.RxEN        =   1'b1;
    uin_hdlc.TxEN        =   1'b1;

    TbErrorCnt = 0;

    #1000ns;
    uin_hdlc.Rst         =   1'b1;
  endtask

  task WriteAddress(input logic [2:0] Address ,input logic [7:0] Data);
    @(posedge uin_hdlc.Clk);
    uin_hdlc.Address     = Address;
    uin_hdlc.WriteEnable = 1'b1;
    uin_hdlc.DataIn      = Data;
    uin_hdlc.Rx          = uin_hdlc.Tx; //Added to keep transfering Tx to Rx during write.
    @(posedge uin_hdlc.Clk);
    uin_hdlc.Rx          = uin_hdlc.Tx; //Added to keep transfering Tx to Rx during write.
    uin_hdlc.WriteEnable = 1'b0;
  endtask

  task ReadAddress(input logic [2:0] Address ,output logic [7:0] Data);
    @(posedge uin_hdlc.Clk);
    uin_hdlc.Address    = Address;
    uin_hdlc.ReadEnable = 1'b1;
    #100ns;
    Data                = uin_hdlc.DataOut;
    @(posedge uin_hdlc.Clk);
    uin_hdlc.ReadEnable = 1'b0;
  endtask


  task Receive();
    logic [7:0] ReadData;

    //RX flag
    @(posedge uin_hdlc.Clk);
    uin_hdlc.Rx = 1'b0;
    @(posedge uin_hdlc.Clk);
    uin_hdlc.Rx = 1'b1;
    @(posedge uin_hdlc.Clk);
    uin_hdlc.Rx = 1'b1;
    @(posedge uin_hdlc.Clk);
    uin_hdlc.Rx = 1'b1;
    @(posedge uin_hdlc.Clk);
    uin_hdlc.Rx = 1'b1;
    @(posedge uin_hdlc.Clk);
    uin_hdlc.Rx = 1'b1;
    @(posedge uin_hdlc.Clk);
    uin_hdlc.Rx = 1'b1;
    @(posedge uin_hdlc.Clk);
    uin_hdlc.Rx = 1'b0;
    @(posedge uin_hdlc.Clk);
    uin_hdlc.Rx = 1'b1;
@(posedge uin_hdlc.Clk);
    uin_hdlc.Address = 1'h2;
@(posedge uin_hdlc.Clk);
    uin_hdlc.Address = 1'h2;

    repeat(8)
      @(posedge uin_hdlc.Clk);

    ReadAddress(3'b010 , ReadData);
    $display("Rx_SC=%h", ReadData);

  endtask
    
  


  task Verification9();
  logic [7:0] writeData;
  logic [7:0] dataIn;
  logic [7:0] transmitData;
  transmitData = 8'b0000000;
  dataIn = 8'b10101010;
  writeData = 8'b00000100;
  for(int i = 0; i < 126; i=i+1) begin
    WriteAddress(TX_BUFF, dataIn);
  end
  WriteAddress(3'b000, transmitData);
  WriteAddress(3'b000, 8'b0000000);
  for(int i = 0; i < 30; i=i+1) begin
      @(posedge uin_hdlc.Clk);
    //#20;
  end
  WriteAddress(3'b000, writeData);
  for(int i = 0; i < 12600; i=i+1) begin
      @(posedge uin_hdlc.Clk);
  end
  @(posedge uin_hdlc.Clk);
  @(posedge uin_hdlc.Clk);
  @(posedge uin_hdlc.Clk);
  @(posedge uin_hdlc.Clk);
  @(posedge uin_hdlc.Clk);
  @(posedge uin_hdlc.Clk);
  endtask

  task Verification17();
    // data_hdlc inputValue;
    logic [7:0] readData;
    logic [7:0] dataIn;
    logic [7:0] transmitData;
    dataIn = 8'b10101010;
    transmitData = 8'b0000010;
    for(int i = 0; i < 126; i=i+1) begin
      WriteAddress(3'b001, dataIn);
      //#20;
		end
    WriteAddress(3'b000, transmitData);
    for(int i = 0; i < 12600; i=i+1) begin
        @(posedge uin_hdlc.Clk);
      //#20;
		end
    @(posedge uin_hdlc.Clk);
    @(posedge uin_hdlc.Clk);
    @(posedge uin_hdlc.Clk);
    ReadAddress(3'b000, readData);
    $display("Tx_SC=%b", readData);

  endtask

  task Verification6();
    // data_hdlc inputValue;
    logic [7:0] readData;
    logic [7:0] dataIn;
    logic [7:0] transmitData;
    dataIn = 255;
    transmitData = 8'b0000010;
    for(int j = 0; j < 40; j=j+1) begin
      //#20;
        ReadAddress(3'b001, readData);
        WriteAddress(3'b001, dataIn);
                uin_hdlc.Rx = uin_hdlc.Tx;
	end
    WriteAddress(3'b001, dataIn);
    
    WriteAddress(3'b000, dataIn);
    repeat(10)
        @(posedge uin_hdlc.Clk)
    for(int j = 0; j < 40; j=j+1) begin
      //#20;
            uin_hdlc.Rx = uin_hdlc.Tx;

	end

    @(posedge uin_hdlc.Clk);
    @(posedge uin_hdlc.Clk);
    @(posedge uin_hdlc.Clk);
    ReadAddress(3'b001, readData);
    $display("Tx_SC=%b", readData);

  endtask

 task Verification8();      //Used for generating increasing data_in and aborting at a certain point in time, if desired.
    // data_hdlc inputValue;
    logic [7:0] readData;
    logic [7:0] dataIn;
    logic [7:0] transmitData;
    logic [7:0] receiveData;
    dataIn = 8'b10101010;
    transmitData = 8'b0000010;
    receiveData = 8'b0000010;
    for(int i = 0; i < 126; i=i+1) begin
      WriteAddress(TX_BUFF, 255);                  //Write the data to register 1
		end
    WriteAddress(TX_SC, transmitData);         //Start transfer
    for(int i = 0; i < 2500; i=i+1) begin
       /* if(i==1500) begin
            transmitData = 8'b00000100;
            WriteAddress(3'b000, transmitData);
        end*/
        @(posedge uin_hdlc.Clk);
        uin_hdlc.Rx = uin_hdlc.Tx;
      //#20;
	end
    @(posedge uin_hdlc.Clk);
    @(posedge uin_hdlc.Clk);
    @(posedge uin_hdlc.Clk);
    ReadAddress(RX_SC, readData);
    $display("Rx_SC=%b", readData);

  endtask

  task random_input();
    automatic logic[7:0] Data = '0;
    logic [7:0] size;

    size = $urandom_range(1, 126); 
    //Generate random data and write it to TX_buffer
    for (int i = 0; i < size; i++) begin
        Data = $urandom();
        WriteAddress(TX_BUFF, Data);
    end
    $display("%d bytes of data written to TX_BUFF", size);
    //Initiate transfer
    WriteAddress(TX_SC, TX_ENABLE);  
    for(int i = 0; i < 2200; i=i+1) begin
       /* if(i==1500) begin
            transmitData = 8'b00000100;
            WriteAddress(3'b000, transmitData);
        end*/
        @(posedge uin_hdlc.Clk);
        uin_hdlc.Rx = uin_hdlc.Tx;
      //#20;
	end
    

  endtask


  task Verification1_Error();
    logic [7:0] readData;
    logic [7:0] writeData;

    writeData = 8'b00100000;
    WriteAddress(3'b010, writeData);

  uin_hdlc.Rx = 1'b0;
  @(posedge uin_hdlc.Clk);
  uin_hdlc.Rx = 1'b1;
  @(posedge uin_hdlc.Clk);
  uin_hdlc.Rx = 1'b1;
  @(posedge uin_hdlc.Clk);
  uin_hdlc.Rx = 1'b1;
  @(posedge uin_hdlc.Clk);
  uin_hdlc.Rx = 1'b1;
  @(posedge uin_hdlc.Clk);
  uin_hdlc.Rx = 1'b1;
  @(posedge uin_hdlc.Clk);
  uin_hdlc.Rx = 1'b1;
  @(posedge uin_hdlc.Clk);
  uin_hdlc.Rx = 1'b0;
  @(posedge uin_hdlc.Clk);

uin_hdlc.Rx = 1'b1;
@(posedge uin_hdlc.Clk);
uin_hdlc.Rx = 1'b0;
@(posedge uin_hdlc.Clk);
uin_hdlc.Rx = 1'b1;
@(posedge uin_hdlc.Clk);
uin_hdlc.Rx = 1'b0;
@(posedge uin_hdlc.Clk);
uin_hdlc.Rx = 1'b1;
@(posedge uin_hdlc.Clk);
uin_hdlc.Rx = 1'b0;
@(posedge uin_hdlc.Clk);
uin_hdlc.Rx = 1'b1;
@(posedge uin_hdlc.Clk);
uin_hdlc.Rx = 1'b0;
@(posedge uin_hdlc.Clk);

uin_hdlc.Rx = 1'b0;
@(posedge uin_hdlc.Clk);
uin_hdlc.Rx = 1'b0;
@(posedge uin_hdlc.Clk);
uin_hdlc.Rx = 1'b0;
@(posedge uin_hdlc.Clk);
uin_hdlc.Rx = 1'b0;
@(posedge uin_hdlc.Clk);
uin_hdlc.Rx = 1'b0;
@(posedge uin_hdlc.Clk);
uin_hdlc.Rx = 1'b0;
@(posedge uin_hdlc.Clk);
uin_hdlc.Rx = 1'b0;
@(posedge uin_hdlc.Clk);
uin_hdlc.Rx = 1'b1;
@(posedge uin_hdlc.Clk);

uin_hdlc.Rx = 1'b1;
@(posedge uin_hdlc.Clk);
uin_hdlc.Rx = 1'b0;
@(posedge uin_hdlc.Clk);
uin_hdlc.Rx = 1'b1;
@(posedge uin_hdlc.Clk);
uin_hdlc.Rx = 1'b0;
@(posedge uin_hdlc.Clk);
uin_hdlc.Rx = 1'b1;
@(posedge uin_hdlc.Clk);
uin_hdlc.Rx = 1'b0;
@(posedge uin_hdlc.Clk);
uin_hdlc.Rx = 1'b1;
@(posedge uin_hdlc.Clk);
uin_hdlc.Rx = 1'b0;
@(posedge uin_hdlc.Clk);


// uin_hdlc.Rx = 1'b1;
// @(posedge uin_hdlc.Clk);
// uin_hdlc.Rx = 1'b1;
// @(posedge uin_hdlc.Clk);
// uin_hdlc.Rx = 1'b1;
// @(posedge uin_hdlc.Clk);
// uin_hdlc.Rx = 1'b1;
// @(posedge uin_hdlc.Clk);
// uin_hdlc.Rx = 1'b0;
// @(posedge uin_hdlc.Clk);
// uin_hdlc.Rx = 1'b0;
// @(posedge uin_hdlc.Clk);
// uin_hdlc.Rx = 1'b0;
// @(posedge uin_hdlc.Clk);
// uin_hdlc.Rx = 1'b0;
// @(posedge uin_hdlc.Clk);
// uin_hdlc.Rx = 1'b0;
// @(posedge uin_hdlc.Clk);
// uin_hdlc.Rx = 1'b0;
// @(posedge uin_hdlc.Clk);
// uin_hdlc.Rx = 1'b0;
// @(posedge uin_hdlc.Clk);
// uin_hdlc.Rx = 1'b0;
// @(posedge uin_hdlc.Clk);
// uin_hdlc.Rx = 1'b1;
// @(posedge uin_hdlc.Clk);
// uin_hdlc.Rx = 1'b1;
// @(posedge uin_hdlc.Clk);
// uin_hdlc.Rx = 1'b1;
// @(posedge uin_hdlc.Clk);
// uin_hdlc.Rx = 1'b1;
// @(posedge uin_hdlc.Clk);

// uin_hdlc.Rx = 1'b0;
// @(posedge uin_hdlc.Clk);
// uin_hdlc.Rx = 1'b0;
// @(posedge uin_hdlc.Clk);
// uin_hdlc.Rx = 1'b0;
// @(posedge uin_hdlc.Clk);
// uin_hdlc.Rx = 1'b0;
// @(posedge uin_hdlc.Clk);
// uin_hdlc.Rx = 1'b0;
// @(posedge uin_hdlc.Clk);
// uin_hdlc.Rx = 1'b0;
// @(posedge uin_hdlc.Clk);
// uin_hdlc.Rx = 1'b0;
// @(posedge uin_hdlc.Clk);
// uin_hdlc.Rx = 1'b0;
// @(posedge uin_hdlc.Clk);
// uin_hdlc.Rx = 1'b0;
// @(posedge uin_hdlc.Clk);
// uin_hdlc.Rx = 1'b0;
// @(posedge uin_hdlc.Clk);
// uin_hdlc.Rx = 1'b0;
// @(posedge uin_hdlc.Clk);
// uin_hdlc.Rx = 1'b0;
// @(posedge uin_hdlc.Clk);
// uin_hdlc.Rx = 1'b0;
// @(posedge uin_hdlc.Clk);
// uin_hdlc.Rx = 1'b0;
// @(posedge uin_hdlc.Clk);
// uin_hdlc.Rx = 1'b0;
// @(posedge uin_hdlc.Clk);
// uin_hdlc.Rx = 1'b0;
// @(posedge uin_hdlc.Clk);

//CRC Code
uin_hdlc.Rx = 1'b0;
@(posedge uin_hdlc.Clk);
uin_hdlc.Rx = 1'b0;
@(posedge uin_hdlc.Clk);
uin_hdlc.Rx = 1'b0;
@(posedge uin_hdlc.Clk);
uin_hdlc.Rx = 1'b0;
@(posedge uin_hdlc.Clk);
uin_hdlc.Rx = 1'b0;
@(posedge uin_hdlc.Clk);
uin_hdlc.Rx = 1'b0;
@(posedge uin_hdlc.Clk);
uin_hdlc.Rx = 1'b0;
@(posedge uin_hdlc.Clk);
uin_hdlc.Rx = 1'b0;
@(posedge uin_hdlc.Clk);
uin_hdlc.Rx = 1'b1;
@(posedge uin_hdlc.Clk);
uin_hdlc.Rx = 1'b0;
@(posedge uin_hdlc.Clk);
uin_hdlc.Rx = 1'b1;
@(posedge uin_hdlc.Clk);
uin_hdlc.Rx = 1'b0;
@(posedge uin_hdlc.Clk);
uin_hdlc.Rx = 1'b1;
@(posedge uin_hdlc.Clk);
uin_hdlc.Rx = 1'b0;
@(posedge uin_hdlc.Clk);
uin_hdlc.Rx = 1'b1;
@(posedge uin_hdlc.Clk);
uin_hdlc.Rx = 1'b0;
@(posedge uin_hdlc.Clk);


uin_hdlc.Rx = 1'b0;
@(posedge uin_hdlc.Clk);
uin_hdlc.Rx = 1'b1;
@(posedge uin_hdlc.Clk);
uin_hdlc.Rx = 1'b1;
@(posedge uin_hdlc.Clk);
uin_hdlc.Rx = 1'b1;
@(posedge uin_hdlc.Clk);
uin_hdlc.Rx = 1'b1;
@(posedge uin_hdlc.Clk);
uin_hdlc.Rx = 1'b1;
@(posedge uin_hdlc.Clk);
uin_hdlc.Rx = 1'b1;
@(posedge uin_hdlc.Clk);
uin_hdlc.Rx = 1'b0;
@(posedge uin_hdlc.Clk);
uin_hdlc.Rx = 1'b1;
//ABORT FRAME
// uin_hdlc.Rx = 1'b1;
// @(posedge uin_hdlc.Clk);
// uin_hdlc.Rx = 1'b1;
// @(posedge uin_hdlc.Clk);
// uin_hdlc.Rx = 1'b1;
// @(posedge uin_hdlc.Clk);
// uin_hdlc.Rx = 1'b1;
// @(posedge uin_hdlc.Clk);
// uin_hdlc.Rx = 1'b1;
// @(posedge uin_hdlc.Clk);
// uin_hdlc.Rx = 1'b1;
// @(posedge uin_hdlc.Clk);
// uin_hdlc.Rx = 1'b1;
// @(posedge uin_hdlc.Clk);
// uin_hdlc.Rx = 1'b0;
// @(posedge uin_hdlc.Clk);

  ReadAddress(3'b011, readData);
  $display("Rx_SC=%b", readData);
  ReadAddress(3'b011, readData);
  $display("Rx_SC=%b", readData);
  ReadAddress(3'b011, readData);
  $display("Rx_SC=%b", readData);
  ReadAddress(3'b011, readData);
  $display("Rx_SC=%b", readData);
  ReadAddress(3'b011, readData);
  $display("Rx_SC=%b", readData);
  ReadAddress(3'b011, readData);
  $display("Rx_SC=%b", readData);
  ReadAddress(3'b011, readData);
  $display("Rx_SC=%b", readData);
  ReadAddress(3'b011, readData);
  $display("Rx_SC=%b", readData);
  ReadAddress(3'b011, readData);
  $display("Rx_SC=%b", readData);
  ReadAddress(3'b011, readData);
  $display("Rx_SC=%b", readData);
  @(posedge uin_hdlc.Clk);
  @(posedge uin_hdlc.Clk);
  @(posedge uin_hdlc.Clk);
  @(posedge uin_hdlc.Clk);
  @(posedge uin_hdlc.Clk);
  @(posedge uin_hdlc.Clk);
  @(posedge uin_hdlc.Clk);
  ReadAddress(3'b011, readData);
  $display("Rx_Data=%b", readData);
  endtask


  task Verification1_Drop();


    logic [7:0] readData;
    logic [7:0] writeData;

  uin_hdlc.Rx = 1'b0;
  @(posedge uin_hdlc.Clk);
  uin_hdlc.Rx = 1'b1;
  @(posedge uin_hdlc.Clk);
  uin_hdlc.Rx = 1'b1;
  @(posedge uin_hdlc.Clk);
  uin_hdlc.Rx = 1'b1;
  @(posedge uin_hdlc.Clk);
  uin_hdlc.Rx = 1'b1;
  @(posedge uin_hdlc.Clk);
  uin_hdlc.Rx = 1'b1;
  @(posedge uin_hdlc.Clk);
  uin_hdlc.Rx = 1'b1;
  @(posedge uin_hdlc.Clk);
  uin_hdlc.Rx = 1'b0;
  @(posedge uin_hdlc.Clk);

uin_hdlc.Rx = 1'b1;
@(posedge uin_hdlc.Clk);
uin_hdlc.Rx = 1'b0;
@(posedge uin_hdlc.Clk);
uin_hdlc.Rx = 1'b1;
@(posedge uin_hdlc.Clk);
uin_hdlc.Rx = 1'b0;
@(posedge uin_hdlc.Clk);
uin_hdlc.Rx = 1'b1;
@(posedge uin_hdlc.Clk);
uin_hdlc.Rx = 1'b0;
@(posedge uin_hdlc.Clk);
uin_hdlc.Rx = 1'b1;
@(posedge uin_hdlc.Clk);
uin_hdlc.Rx = 1'b0;
@(posedge uin_hdlc.Clk);

uin_hdlc.Rx = 1'b0;
@(posedge uin_hdlc.Clk);
uin_hdlc.Rx = 1'b0;
@(posedge uin_hdlc.Clk);
uin_hdlc.Rx = 1'b0;
@(posedge uin_hdlc.Clk);
uin_hdlc.Rx = 1'b0;
@(posedge uin_hdlc.Clk);
uin_hdlc.Rx = 1'b0;
@(posedge uin_hdlc.Clk);
uin_hdlc.Rx = 1'b0;
@(posedge uin_hdlc.Clk);
uin_hdlc.Rx = 1'b0;
@(posedge uin_hdlc.Clk);
uin_hdlc.Rx = 1'b1;
@(posedge uin_hdlc.Clk);

uin_hdlc.Rx = 1'b1;
@(posedge uin_hdlc.Clk);
uin_hdlc.Rx = 1'b0;
@(posedge uin_hdlc.Clk);
uin_hdlc.Rx = 1'b1;
@(posedge uin_hdlc.Clk);
uin_hdlc.Rx = 1'b0;
@(posedge uin_hdlc.Clk);
uin_hdlc.Rx = 1'b1;
@(posedge uin_hdlc.Clk);
uin_hdlc.Rx = 1'b0;
@(posedge uin_hdlc.Clk);
uin_hdlc.Rx = 1'b1;
@(posedge uin_hdlc.Clk);
uin_hdlc.Rx = 1'b0;
@(posedge uin_hdlc.Clk);


uin_hdlc.Rx = 1'b1;
@(posedge uin_hdlc.Clk);
uin_hdlc.Rx = 1'b1;
@(posedge uin_hdlc.Clk);
uin_hdlc.Rx = 1'b1;
@(posedge uin_hdlc.Clk);
uin_hdlc.Rx = 1'b1;
@(posedge uin_hdlc.Clk);
uin_hdlc.Rx = 1'b0;
@(posedge uin_hdlc.Clk);
uin_hdlc.Rx = 1'b0;
@(posedge uin_hdlc.Clk);
uin_hdlc.Rx = 1'b0;
@(posedge uin_hdlc.Clk);
uin_hdlc.Rx = 1'b0;
@(posedge uin_hdlc.Clk);
uin_hdlc.Rx = 1'b0;
@(posedge uin_hdlc.Clk);
uin_hdlc.Rx = 1'b0;
@(posedge uin_hdlc.Clk);
uin_hdlc.Rx = 1'b0;
@(posedge uin_hdlc.Clk);
uin_hdlc.Rx = 1'b0;
@(posedge uin_hdlc.Clk);
uin_hdlc.Rx = 1'b1;
@(posedge uin_hdlc.Clk);
uin_hdlc.Rx = 1'b1;
@(posedge uin_hdlc.Clk);
uin_hdlc.Rx = 1'b1;
@(posedge uin_hdlc.Clk);
uin_hdlc.Rx = 1'b1;
@(posedge uin_hdlc.Clk);

uin_hdlc.Rx = 1'b0;
@(posedge uin_hdlc.Clk);
uin_hdlc.Rx = 1'b1;
@(posedge uin_hdlc.Clk);
uin_hdlc.Rx = 1'b1;
@(posedge uin_hdlc.Clk);
uin_hdlc.Rx = 1'b1;
@(posedge uin_hdlc.Clk);
uin_hdlc.Rx = 1'b1;
@(posedge uin_hdlc.Clk);
uin_hdlc.Rx = 1'b1;
@(posedge uin_hdlc.Clk);
uin_hdlc.Rx = 1'b1;
@(posedge uin_hdlc.Clk);
uin_hdlc.Rx = 1'b0;
@(posedge uin_hdlc.Clk);

//ABORT FRAME
// uin_hdlc.Rx = 1'b1;
// @(posedge uin_hdlc.Clk);
// uin_hdlc.Rx = 1'b1;
// @(posedge uin_hdlc.Clk);
// uin_hdlc.Rx = 1'b1;
// @(posedge uin_hdlc.Clk);
// uin_hdlc.Rx = 1'b1;
// @(posedge uin_hdlc.Clk);
// uin_hdlc.Rx = 1'b1;
// @(posedge uin_hdlc.Clk);
// uin_hdlc.Rx = 1'b1;
// @(posedge uin_hdlc.Clk);
// uin_hdlc.Rx = 1'b1;
// @(posedge uin_hdlc.Clk);
// uin_hdlc.Rx = 1'b0;
// @(posedge uin_hdlc.Clk);


  writeData = 8'b00000000;
  WriteAddress(3'b010, writeData);
  ReadAddress(3'b010, readData);
  $display("Rx_SC=%b", readData);
  @(posedge uin_hdlc.Clk);
  @(posedge uin_hdlc.Clk);
  @(posedge uin_hdlc.Clk);
  @(posedge uin_hdlc.Clk);
  @(posedge uin_hdlc.Clk);
  @(posedge uin_hdlc.Clk);


  uin_hdlc.Address     = 3'b010;
  uin_hdlc.WriteEnable = 1'b1;
  uin_hdlc.DataIn      = 8'b00000010;
  @(posedge uin_hdlc.Clk);
  ReadAddress(3'b011, readData);
  $display("Rx_Data=%b", readData);
  endtask


  task Verification1_Abort();


    logic [7:0] readData;
    logic [7:0] writeData;

  uin_hdlc.Rx = 1'b0;
  @(posedge uin_hdlc.Clk);
  uin_hdlc.Rx = 1'b1;
  @(posedge uin_hdlc.Clk);
  uin_hdlc.Rx = 1'b1;
  @(posedge uin_hdlc.Clk);
  uin_hdlc.Rx = 1'b1;
  @(posedge uin_hdlc.Clk);
  uin_hdlc.Rx = 1'b1;
  @(posedge uin_hdlc.Clk);
  uin_hdlc.Rx = 1'b1;
  @(posedge uin_hdlc.Clk);
  uin_hdlc.Rx = 1'b1;
  @(posedge uin_hdlc.Clk);
  uin_hdlc.Rx = 1'b0;
  @(posedge uin_hdlc.Clk);

uin_hdlc.Rx = 1'b1;
@(posedge uin_hdlc.Clk);
uin_hdlc.Rx = 1'b0;
@(posedge uin_hdlc.Clk);
uin_hdlc.Rx = 1'b1;
@(posedge uin_hdlc.Clk);
uin_hdlc.Rx = 1'b0;
@(posedge uin_hdlc.Clk);
uin_hdlc.Rx = 1'b1;
@(posedge uin_hdlc.Clk);
uin_hdlc.Rx = 1'b0;
@(posedge uin_hdlc.Clk);
uin_hdlc.Rx = 1'b1;
@(posedge uin_hdlc.Clk);
uin_hdlc.Rx = 1'b0;
@(posedge uin_hdlc.Clk);

uin_hdlc.Rx = 1'b0;
@(posedge uin_hdlc.Clk);
uin_hdlc.Rx = 1'b0;
@(posedge uin_hdlc.Clk);
uin_hdlc.Rx = 1'b0;
@(posedge uin_hdlc.Clk);
uin_hdlc.Rx = 1'b0;
@(posedge uin_hdlc.Clk);
uin_hdlc.Rx = 1'b0;
@(posedge uin_hdlc.Clk);
uin_hdlc.Rx = 1'b0;
@(posedge uin_hdlc.Clk);
uin_hdlc.Rx = 1'b0;
@(posedge uin_hdlc.Clk);
uin_hdlc.Rx = 1'b1;
@(posedge uin_hdlc.Clk);

uin_hdlc.Rx = 1'b1;
@(posedge uin_hdlc.Clk);
uin_hdlc.Rx = 1'b0;
@(posedge uin_hdlc.Clk);
uin_hdlc.Rx = 1'b1;
@(posedge uin_hdlc.Clk);
uin_hdlc.Rx = 1'b0;
@(posedge uin_hdlc.Clk);
uin_hdlc.Rx = 1'b1;
@(posedge uin_hdlc.Clk);
uin_hdlc.Rx = 1'b0;
@(posedge uin_hdlc.Clk);
uin_hdlc.Rx = 1'b1;
@(posedge uin_hdlc.Clk);
uin_hdlc.Rx = 1'b0;
@(posedge uin_hdlc.Clk);


uin_hdlc.Rx = 1'b1;
@(posedge uin_hdlc.Clk);
uin_hdlc.Rx = 1'b1;
@(posedge uin_hdlc.Clk);
uin_hdlc.Rx = 1'b1;
@(posedge uin_hdlc.Clk);
uin_hdlc.Rx = 1'b1;
@(posedge uin_hdlc.Clk);
uin_hdlc.Rx = 1'b0;
@(posedge uin_hdlc.Clk);
uin_hdlc.Rx = 1'b0;
@(posedge uin_hdlc.Clk);
uin_hdlc.Rx = 1'b0;
@(posedge uin_hdlc.Clk);
uin_hdlc.Rx = 1'b0;
@(posedge uin_hdlc.Clk);
uin_hdlc.Rx = 1'b0;
@(posedge uin_hdlc.Clk);
uin_hdlc.Rx = 1'b0;
@(posedge uin_hdlc.Clk);
uin_hdlc.Rx = 1'b0;
@(posedge uin_hdlc.Clk);
uin_hdlc.Rx = 1'b0;
@(posedge uin_hdlc.Clk);
uin_hdlc.Rx = 1'b1;
@(posedge uin_hdlc.Clk);
uin_hdlc.Rx = 1'b1;
@(posedge uin_hdlc.Clk);
uin_hdlc.Rx = 1'b1;
@(posedge uin_hdlc.Clk);
uin_hdlc.Rx = 1'b1;
@(posedge uin_hdlc.Clk);

// uin_hdlc.Rx = 1'b0;
// @(posedge uin_hdlc.Clk);
// uin_hdlc.Rx = 1'b1;
// @(posedge uin_hdlc.Clk);
// uin_hdlc.Rx = 1'b1;
// @(posedge uin_hdlc.Clk);
// uin_hdlc.Rx = 1'b1;
// @(posedge uin_hdlc.Clk);
// uin_hdlc.Rx = 1'b1;
// @(posedge uin_hdlc.Clk);
// uin_hdlc.Rx = 1'b1;
// @(posedge uin_hdlc.Clk);
// uin_hdlc.Rx = 1'b1;
// @(posedge uin_hdlc.Clk);
// uin_hdlc.Rx = 1'b0;
// @(posedge uin_hdlc.Clk);

//ABORT FRAME
uin_hdlc.Rx = 1'b1;
@(posedge uin_hdlc.Clk);
uin_hdlc.Rx = 1'b1;
@(posedge uin_hdlc.Clk);
uin_hdlc.Rx = 1'b1;
@(posedge uin_hdlc.Clk);
uin_hdlc.Rx = 1'b1;
@(posedge uin_hdlc.Clk);
uin_hdlc.Rx = 1'b1;
@(posedge uin_hdlc.Clk);
uin_hdlc.Rx = 1'b1;
@(posedge uin_hdlc.Clk);
uin_hdlc.Rx = 1'b1;
@(posedge uin_hdlc.Clk);
uin_hdlc.Rx = 1'b0;
@(posedge uin_hdlc.Clk);


  @(posedge uin_hdlc.Clk);
  @(posedge uin_hdlc.Clk);
  @(posedge uin_hdlc.Clk);
  @(posedge uin_hdlc.Clk);
  @(posedge uin_hdlc.Clk);
  @(posedge uin_hdlc.Clk);
  @(posedge uin_hdlc.Clk);

  ReadAddress(3'b011, readData);
  $display("Rx_Data=%b", readData);
  endtask

endprogram
